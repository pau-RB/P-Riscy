import Types::*;
import ProcTypes::*;

(* noinline *)
function Data alu(Data a, Data b, AluFunc func);

    Data res = case(func)
        Add   : (a + b);
        Sub   : (a - b);
        And   : (a & b);
        Or    : (a | b);
        Xor   : (a ^ b);
        Slt   : zeroExtend( pack( signedLT(a, b) ) );
        Sltu  : zeroExtend( pack( a < b ) );
        // 5-bit shift width for 32-bit data
        Sll   : (a << b[4:0]);
        Srl   : (a >> b[4:0]);
        Sra   : signedShiftRight(a, b[4:0]);
    endcase;

    return res;

endfunction

(* noinline *)
function Bool aluBr(Data a, Data b, BrFunc brFunc);

    Bool brTaken = case(brFunc)
        Eq  : (a == b);
        Neq : (a != b);
        Lt  : signedLT(a, b);
        Ltu : (a < b);
        Ge  : signedGE(a, b);
        Geu : (a >= b);
        AT  : True;
        NT  : False;
    endcase;

    return brTaken;

endfunction

(* noinline *)
function Addr brAddrCalc(Addr pc, Data val, IType iType, Data imm, Bool taken);

    Addr pcPlus4 = pc + 4;
    Addr targetAddr = case (iType)
        J   : (pc + imm);
        Fork: (pc + imm);
        Jr  : {truncateLSB(val + imm), 1'b0};
        Forkr: {truncateLSB(val + imm), 1'b0};
        Br  : (taken ? pc + imm : pcPlus4);
        default: pcPlus4;
    endcase;

    return targetAddr;

endfunction