import Types::*;
import Memory::*;
import Vector::*;
import ProcTypes::*;
import MemTypes::*;


//////////// LOCAL DATA-BASED MEMORY ////////////

typedef enum{Ld, St}  MemOp  deriving(Eq, Bits, FShow);

typedef struct{
    MemOp     op;
    Addr      addr;
    Data      data;
    StoreFunc func;
} MemReq deriving(Eq, Bits, FShow);

typedef Data MemResp;

interface Cache;
    method Action req(MemReq r);
    method ActionValue#(MemResp) resp;
endinterface