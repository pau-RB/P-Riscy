import Types::*;
import ProcTypes::*;
import MemTypes::*;
import Fifo::*;
import Ehr::*;


typedef Bit#(TSub#(AddrSz,TLog#(CacheLineBytes))) CacheLineNum;

typedef enum {
	Full,
	Evict,
	Ghost,
	Dry,
	Empty
} StreamStatus deriving(Bits, Eq, FShow);


interface Stream;

	// Flow control
	method ActionValue#(DecToken) fetch();
	method Action                 redirect(Redirect r);

	// Thread control
	method Bool                   available();
	method Action                 start(Addr sPC, Addr sFP);
	method Action                 evict();
	method Action                 backendDry();

	// Debug
	method StreamStatus           currentState();
	method Addr                   currentPC();
	method Addr                   currentFP();
	method Addr                   decodePC();
	method Bool                   notEmpty();
	method Bool                   isl0Ihit();

endinterface

// evict < {Redirect, Fetch} < l1I_resp < l1I_req < do_dry < start
// Redirect C Fetch
// Redirect C do_dry
module mkStream (WideMem l1I, Stream ifc);

	Ehr#(3,StreamStatus)   state     <- mkEhr(Empty);
	Ehr#(2,Addr)           pc        <- mkEhr('0);
	Reg#(Addr)             fp        <- mkReg('0);
	Reg#(Bool)             epoch     <- mkReg(False);

	Fifo#(1,DecToken)      inst      <- mkStageFifo();
	Fifo#(1,Redirect)      redirectQ <- mkBypassFifo();
	Fifo#(1,void)          dryQ      <- mkBypassFifo();
	
	Reg #(CacheLine)       l0I       <- mkRegU();
	Reg #(CacheLineNum)    l0Iline   <- mkRegU();
	Reg #(Bool)            l0Ival    <- mkReg(False);
	Fifo#(1, CacheLineNum) l1Ireq    <- mkPipelineFifo();

	// Note: After pc+4 we might request a new line. Then, we might receive
	// a redirect request and generate a new L1I request. When getting the
	// responses, we will only keep the last ones

	CacheLineNum pcline = truncateLSB(pc[0]);
	Bool l0Ihit = (pcline==l0Iline)&&l0Ival;

	// 0 - Interact with L1I

	rule do_l1Ireq;

		CacheLineNum nextpcline = truncateLSB(pc[1]);

		if(nextpcline != l0Iline) begin
    		l1I.req(WideMemReq {
        	        		write_en: '0,
        	        		addr:     {nextpcline,'0},
        	        		data:     ?             });
    		l1Ireq.enq(pcline);
    	end

	endrule

	rule do_l1Iresp;

		CacheLine data <- l1I.resp();

		l0I     <= data;
		l0Iline <= l1Ireq.first(); l1Ireq.deq();
		l0Ival  <= True;

	endrule
	

	// 1 - Consider redirect

	rule do_redirect if (state[1] == Full || state[1] == Evict || state[1] == Ghost || state[1] == Dry);

		// Do redirect
		let redirect = redirectQ.first(); redirectQ.deq();
		pc[0] <= redirect.nextPc;
		epoch <= redirect.epoch;

		if(state[1] == Evict || state[1] == Dry) begin
			state[1] <= Ghost;
		end

	endrule


	// 2 - Try to fetch

	rule do_fetch if ((state[1] == Full && l0Ihit) || state[1] == Evict || state[1] == Ghost);

		if(state[1] == Full && l0Ihit) begin

			// Fetch real instruction
			CacheWordSelect wordSelect = truncate(pc[0] >> 2);
			inst.enq(DecToken{ inst:  l0I[wordSelect],
							   pc:    pc[0],
							   fp:    fp,
							   ghost: False,
							   epoch: epoch});
			pc[0] <= pc[0]+4;

		end else if (state[1] == Evict) begin
			
			if(l0Ihit) begin

				// Fetch real instruction
				CacheWordSelect wordSelect = truncate(pc[0] >> 2);
				inst.enq(DecToken{ inst:  l0I[wordSelect],
								   pc:    pc[0],
								   fp:    fp,
								   ghost: False,
								   epoch: epoch});
				pc[0] <= pc[0]+4;

			end else begin
				
				// Fetch ghost
				state[1] <= Dry;
				inst.enq(DecToken{ inst:  ?,
								   pc:    pc[0],
								   fp:    fp,
								   ghost: True,
								   epoch: epoch});

			end

		end else begin
			
			// Fetch ghost
			state[1] <= Dry;
			inst.enq(DecToken{ inst:  ?,
							   pc:    pc[0],
							   fp:    fp,
							   ghost: True,
							   epoch: epoch});

		end

	endrule

	// 3 - Check if pipeline is flush

	rule do_dry if(state[1] == Dry);

		dryQ.deq();
		state[1] <= Empty;

	endrule

	// 4 - Consider external requests

	method Bool available();
		return (state[2] == Empty);
	endmethod

	method Action start(Addr sPC, Addr sFP) if(state[2] == Empty);
		state [2] <= Full;
		pc[1]     <= sPC;
		fp        <= sFP;
		epoch     <= False;
	endmethod


	method Action evict()         if(state[0] == Full);
		state [0] <= Evict;
	endmethod


	method Action backendDry()    if(state[1] == Dry);
		dryQ.enq(?);
	endmethod


	// Attend backend requests

	method ActionValue#(DecToken) fetch();
		DecToken i = inst.first(); inst.deq();
		return i;
	endmethod	

	method Action redirect(Redirect r);
		redirectQ.enq(r);
	endmethod

	method StreamStatus currentState();
		return state[0];
	endmethod

	method Addr currentPC();
		if(state[0] != Empty) begin
			return pc[0];
		end else begin
			return '0;
		end
	endmethod

	method Addr currentFP();
		if(state[0] != Empty) begin
			return fp;
		end else begin
			return '0;
		end
	endmethod

	method Addr decodePC();
		if(inst.notEmpty()) begin
			return inst.first().pc;
		end else begin
			return '0;
		end
	endmethod

	method Bool notEmpty();
		return  inst.notEmpty();
	endmethod

	method Bool isl0Ihit();
		return  l0Ihit;
	endmethod

endmodule