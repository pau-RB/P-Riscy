import Types::*;

// Connectal (FPGA)
Bool wb_ext_DEBUG  = False;
Bool msg_ext_DEBUG = True;

// Verilog (SIM)
Bool msg_DEBUG     = False;
Bool perf_DEBUG    = False;

// MSG relay
typedef  80 THQ_LEN;
Addr     msg_ADDR  = 'h0fff0;
Addr     max_ADDR  = 'h3fffc;

// Main Token Queue
typedef 16 MTQ_LEN;

// Core width
typedef 4 FrontWidth;
typedef Bit#(TLog#(FrontWidth)) FrontID;

// Verification
typedef Bit#(32) VerifID;