`define ConnectalVersion 22.05.23b
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 20
`define DerivedClockPeriod 10.000000
`define CnocTop 
`define XsimHostInterface 
`define PhysAddrWidth 40
`define SIMULATION 
`define SVDPI 
`define CONNECTAL_BITS_DEPENDENCES vlsim
`define BOARD_verilator 
