typedef	1024 CMRTHQ_LEN;